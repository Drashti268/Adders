`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:59:25 05/15/2023 
// Design Name: 
// Module Name:    half_adder_st 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module half_adder_st(a,b,sum,carry);
input a,b;
output sum,carry;
xor x1(sum,a,b);
and a1(carry,a,b);


endmodule
